package designparameters;

parameter SLAVE_SIZE=8;
parameter SLAVE_ADDR=7'b1001100;

endpackage